module top_module (
    output out);
    //assign Gnd=1'b0;
    assign out=1'b0;

endmodule
